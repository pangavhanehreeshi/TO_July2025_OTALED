** sch_path: /foss/designs/thesis/TO_July2025_OTALED/OTALED/design_data/xschem/FMD_QNC_foldedcascode.sch
**.subckt FMD_QNC_foldedcascode AVDD IBIAS PLUS MINUS VOUT AVSS
*.ipin PLUS
*.ipin MINUS
*.ipin AVSS
*.ipin IBIAS
*.ipin AVDD
*.opin VOUT
XM1 net6 MINUS net1 AVDD sg13_lv_pmos w=20u l=2u ng=4 m=1
XM5 net7 net8 net4 AVSS sg13_lv_nmos w=2u l=2u ng=2 m=1
XM2 net4 PLUS net1 AVDD sg13_lv_pmos w=20u l=2u ng=4 m=1
XM3 net2 net7 AVDD AVDD sg13_lv_pmos w=13u l=2u ng=2 m=1
XM4 net3 net7 AVDD AVDD sg13_lv_pmos w=13u l=2u ng=2 m=1
XM7 net7 net9 net2 AVDD sg13_lv_pmos w=8u l=2u ng=4 m=1
XM8 VOUT net9 net3 AVDD sg13_lv_pmos w=8u l=2u ng=4 m=1
XM6 VOUT net8 net6 AVSS sg13_lv_nmos w=2u l=2u ng=2 m=1
XM9 net4 net5 AVSS AVSS sg13_lv_nmos w=4u l=2u ng=2 m=1
XM0 net6 net5 AVSS AVSS sg13_lv_nmos w=4u l=2u ng=2 m=1
XMt net1 net10 AVDD AVDD sg13_lv_pmos w=32u l=5u ng=4 m=1
XM13 IBIAS net7 net5 AVSS sg13_lv_nmos w=4u l=2u ng=2 m=1
XM15 net5 net5 AVSS AVSS sg13_lv_nmos w=4u l=2u ng=1 m=1
XM16 net8 net5 AVSS AVSS sg13_lv_nmos w=4u l=2u ng=1 m=1
XM14 AVDD net7 net8 AVSS sg13_lv_nmos w=15u l=0.5u ng=2 m=1
XM12 net9 net8 AVSS AVSS sg13_lv_nmos w=2u l=2u ng=1 m=1
XM10 net9 net9 AVDD AVDD sg13_lv_pmos w=8u l=2u ng=2 m=1
XM11 net10 net5 AVSS AVSS sg13_lv_nmos w=4u l=2u ng=1 m=1
XMtb net10 net10 AVDD AVDD sg13_lv_pmos w=28u l=5u ng=4 m=1
XM18 net5 AVSS AVSS AVSS sg13_lv_nmos w=4u l=2u ng=1 m=1
XM19 AVDD AVSS AVSS AVSS sg13_lv_nmos w=15u l=0.5u ng=2 m=1
XM20 net4 AVSS AVSS AVSS sg13_lv_nmos w=4u l=2u ng=2 m=1
XM21 net7 AVSS AVSS AVSS sg13_lv_nmos w=2u l=2u ng=2 m=1
XM22 VOUT AVSS AVSS AVSS sg13_lv_nmos w=2u l=2u ng=2 m=1
XM23 AVDD AVDD net1 AVDD sg13_lv_pmos w=10u l=2u ng=2 m=1
XM24 AVDD AVDD net1 AVDD sg13_lv_pmos w=10u l=2u ng=2 m=1
XM25 net10 AVSS AVSS AVSS sg13_lv_nmos w=8u l=2u ng=2 m=1
XM26 net9 AVSS AVSS AVSS sg13_lv_nmos w=4u l=2u ng=2 m=1
XMtb1 net10 AVDD AVDD AVDD sg13_lv_pmos w=14u l=5u ng=2 m=1
XM27 net9 AVDD AVDD AVDD sg13_lv_pmos w=8u l=2u ng=2 m=1
XMt1 net1 AVDD AVDD AVDD sg13_lv_pmos w=16u l=5u ng=2 m=1
XD3 AVDD AVDD AVSS diodevdd_2kv m=1
XD4 AVDD AVDD AVSS diodevss_2kv m=1
XD5 AVDD AVSS AVSS diodevdd_2kv m=1
XD6 AVDD AVSS AVSS diodevss_2kv m=1
XX2 AVSS bondpad size=80u shape=0 padtype=0
XX3 AVDD bondpad size=80u shape=0 padtype=0
XD7 AVDD IBIAS AVSS diodevdd_2kv m=1
XD8 AVDD IBIAS AVSS diodevss_2kv m=1
XX4 IBIAS bondpad size=80u shape=0 padtype=0
XC2 VOUT AVSS cap_cmim w=25.82e-6 l=25.82e-6 m=1
XX1 VOUT bondpad size=80u shape=0 padtype=0
XX5 PLUS bondpad size=80u shape=0 padtype=0
XX6 MINUS bondpad size=80u shape=0 padtype=0
XM30 net8 AVSS AVSS AVSS sg13_lv_nmos w=4u l=2u ng=1 m=1
**.ends
.end
